module Mux2x1_5bits(input [4:0]A,input [4:0] B,input S, output [4:0]Y);
   assign Y = (S==0) ? A:B;
endmodule